library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

   
package my_font is

	Type font_sign_type	is ARRAY (0 to 15) of STD_logic_vector(0 to 15);
	Type font_table_type is ARRAY (0 to 15) of font_sign_type;		 
	
	constant font_table : font_table_type := 
	(
		(		
		"0000000000000000",
		"0000000000000000",
		"0000111111110000",
		"0001111111111000",
		"0001111001111000",
		"0001110000111000",
		"0001110000111000",
		"0001110000111000",
		"0001110000111000",
		"0001110000111000",
		"0001110000111000",
		"0001110000111000",
		"0001111001111000",
		"0001111111111000",
		"0000111111110000",
		"0000000000000000"
		), 
		(		
		"0000000000000000",	
		"0000000000000000",
		"0000000111000000",
		"0000011111000000",
		"0000011111000000",
		"0000000111000000",
		"0000000111000000",
		"0000000111000000",
		"0000000111000000",	
		"0000000111000000",
		"0000000111000000",
		"0000000111000000",
		"0000000111000000",
		"0000111111111000",
		"0000111111111000",
		"0000000000000000"
		), 
		(		
		"0000000000000000",	
		"0000000000000000",
		"0000001111100000",
		"0000011111110000",
		"0000111000111000",
		"0000110000111000",
		"0000000000111000",
		"0000000001110000",
		"0000000011100000",	
		"0000000111000000",
		"0000001110000000",
		"0000011100000000",
		"0000111000000000",
		"0001111111111000",
		"0001111111111000",
		"0000000000000000"
		),
		(		
		"0000000000000000",	
		"0000000000000000",
		"0000011111110000",
		"0000111111111000",
		"0001111000111100",
		"0001110000011100",
		"0000000000011100",
		"0000000000111000",
		"0000000000111000",	
		"0000000000111000",
		"0000000000011100",
		"0001110000011100",
		"0001111000111100",
		"0000111111111000",
		"0000011111110000",
		"0000000000000000"
		), 
		(		
		"0000000000000000",	
		"0000000000000000",
		"0000000011100000",
		"0000000111100000",
		"0000001111100000",
		"0000011101100000",
		"0000111001100000",
		"0001110001100000",
		"0001111111111000",	
		"0000111111110000",
		"0000000001100000",
		"0000000001100000",
		"0000000001100000",
		"0000000001100000",
		"0000000001100000",
		"0000000000000000"
		),
		(		
		"0000000000000000",	
		"0000000000000000",
		"0001111111110000",
		"0001111111110000",
		"0001110000000000",
		"0001110000000000",
		"0001111111000000",
		"0001111111100000",
		"0000000001110000",	
		"0000000000111000",
		"0000000000111000",
		"0001110000111000",
		"0001110000111000",
		"0000111111110000",
		"0000011111100000",
		"0000000000000000"
		), 
		(		
        "0000000000000000",    
        "0000000000000000",
        "0000000011110000",
        "0000001111110000",
        "0000011100000000",
        "0000111000000000",
        "0001110000000000",
        "0001110000000000",
        "0001111111100000",    
        "0001111111110000",
        "0001110000110000",
        "0001110000110000",
        "0001110000110000",
        "0000111111100000",
        "0000011111000000",
        "0000000000000000"
        ), 
		(		
		"0000000000000000",	
		"0000000000000000",
		"0000111111110000",
		"0000111111110000",
		"0000000000110000",
		"0000000001110000",
		"0000000011100000",
		"0000000111000000",
		"0000001110000000",	
		"0000001110000000",
		"0000001100000000",
		"0000001100000000",
		"0000001100000000",
		"0000001100000000",
		"0000001100000000",
		"0000000000000000"
		), 
		(		
        "0000000000000000",    
        "0000000000000000",
        "0000011111100000",
        "0000111111110000",
        "0001111001111000",
        "0001110000111000",
        "0001111001111000",
        "0000111111110000",
        "0000011111100000",    
        "0000111111110000",
        "0001111001111000",
        "0001110000111000",
        "0001111001111000",
        "0000111111110000",
        "0000011111100000",
        "0000000000000000"
        ), 
		(		
        "0000000000000000",
        "0000000000000000", 
        "0000011111000000",
        "0000111111100000",
        "0000110000110000", 
        "0000110000110000",
        "0000110000110000",
        "0000111111110000",
        "0000011111110000", 
        "0000000000110000",  
        "0000000000110000",
        "0000000000110000",
        "0000000011100000",
        "0000111111000000",
        "0000111110000000",           
        "0000000000000000"
        ), 
		(                 --10		
		"0000000000000000",	
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",	
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000011100000",
		"0000000011100000",
		"0000000011100000",
		"0000000000000000"
		),
		(		           --11 
		"0000000000000000",	
		"0000000000000000",
		"0001100000011000",
		"0001100000011000",
		"0001100000011000",
		"0001100000011000",
		"0001100000011000",
		"0001111111111000",
		"0001111111111000",	
		"0001100000011000",
		"0001100000011000",
		"0001100000011000",
		"0001100000011000",
		"0001100000011000",
		"0001100000011000",
		"0000000000000000"
		),
		(		           --12
		"0000000000000000",	
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000111111110000",
		"0000111111110000",	
		"0000000011100000",
		"0000000111000000",
		"0000001110000000",
		"0000011100000000",
		"0000111111110000",
		"0000111111110000",
		"0000000000000000"
		), 
		(		           --13
		"0000000000000000",	
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"1111111111111111",
		"1111111111111111",	
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000"
		),
		(		           --14
		"0000000110000000",	
		"0000000110000000",
		"0000000110000000",
		"0000000110000000",
		"0000000110000000",
		"0000000110000000",
		"0000000110000000",
		"0000000110000000",
		"0000000110000000",	
		"0000000110000000",
		"0000000110000000",
		"0000000110000000",
		"0000000110000000",
		"0000000110000000",
		"0000000110000000",
		"0000000110000000"
		),
		(		           --15
		"0000000000000000",	
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",	
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000"
		)
	);
	
	
end my_font;